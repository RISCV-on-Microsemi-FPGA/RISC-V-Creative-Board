`timescale 1ns/1ns
// ********************************************************************/ 
// Microsemi Corporation Proprietary and Confidential
// Copyright 2014 Microsemi Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED 
// IN ADVANCE IN WRITING.  
//  
//
// CoreSPI User Testbench
//
//
// SVN Revision Information:
// SVN $Revision: 23762 $
// SVN $Date: 2014-11-11 08:01:54 -0800 (Tue, 11 Nov 2014) $
//
// Resolved SARs
// SAR      Date     Who   Description
//
//
// *********************************************************************/ 
module testbench();

`include "../../../../coreparameters.v"

reg  SYSCLK;      
reg  SYSRSTN;     
wire PCLK;        
wire PRESETN;     
wire [31:0] PADDR;      
wire PENABLE;     
wire PWRITE;      
wire [31:0] PWDATA;     
wire [31:0] PRDATA;     
wire [31:0] PRDATA_0;     
wire [31:0] PRDATA_1;     
wire [15:0] PSEL;
         
wire [255:0] INTERRUPT;   
wire [31:0]  GP_OUT;      
wire [31:0]  GP_IN;       
wire FINISHED;  
wire FAILED;

wire Logic0 = 1'b0;
wire Logic1 = 1'b1;    


// ********************************************************************************
// Clocks and Reset


initial
 begin
  SYSRSTN <= 1'b0;
  #100;
  SYSRSTN <= 1'b1;
 end

// Clock is 100MHz
always
 begin
   SYSCLK <= 1'b0;
   #5;
   SYSCLK <= 1'b1;
   #5;
 end

initial
begin
 	// wait until all BFM's are finished
	wait(FINISHED === 1'b1);
	$stop;
	$finish;
end
 
   
// ********************************************************************************
// APB Master  

CORESPI_BFM_APB  #(.VECTFILE     ("user_tb.vec") )
     UBFM (.SYSCLK       (SYSCLK), 
           .SYSRSTN      (SYSRSTN), 
           .PCLK         (PCLK), 
           .PRESETN      (PRESETN), 
           .PADDR        (PADDR), 
           .PENABLE      (PENABLE), 
           .PWRITE       (PWRITE), 
           .PWDATA       (PWDATA), 
           .PRDATA       (PRDATA), 
           .PREADY       (Logic1), 
           .PSLVERR      (Logic0), 
           .PSEL         (PSEL), 
           .INTERRUPT    (INTERRUPT),
           .GP_OUT       (GP_OUT), 
           .GP_IN        (GP_IN), 
           .EXT_WR       (), 
           .EXT_RD       (), 
           .EXT_ADDR     (), 
           .EXT_DATA     (), 
           .EXT_WAIT     (Logic0), 
           .CON_ADDR     (), 
           .CON_DATA     (), 
           .CON_RD       (Logic0), 
           .CON_WR       (Logic0), 
           .CON_BUSY     (), 
           .FINISHED     (FINISHED), 
           .FAILED       (FAILED)
        );                       
                   
assign PRDATA = ( PSEL[1] ? PRDATA_1 : PRDATA_0) ;                   
                         
                         
/* #############################################################################
                         
SPIINT      Output interrupt 
SPISDO      Output serial data out (generated by SPI as master)
SPISS[7:0]  Output slave select (generated by SPI as master)
SPISCLKO    Output shift clock out (generated by SPI as master)
SPISDI      Input  shift data in (master or slave)
SPIRXAVAIL  Output request for data to be read - rx data available
SPITXRFM    Output indicates transmit done - ready for more
SPISSI      Input  slave select (when SPI in slave mode)
SPIOEN      Output output enable (when de-asserted output pad for SPISDO tri-stated). This is active when the SPI is writing output data and deactivated when there is not data to write. This signal is active high.
SPIMode     Output mode:  (when 1,  SPI is master, when 0, SPI is slave)

*/

// ********************************************************************************
// SPI Core - Master    

wire [7:0] M_SPISS;

CORESPI # (
  //.FAMILY              (FAMILY),
  .APB_DWIDTH          (32),
  .CFG_FRAME_SIZE      (32),
  .CFG_FIFO_DEPTH      (4),
  .CFG_CLK             (3),
  .CFG_MODE            (0),
  .CFG_MOT_MODE        (0),
  .CFG_MOT_SSEL        (0),
  .CFG_TI_NSC_CUSTOM   (0),
  .CFG_TI_NSC_FRC      (0),
  .CFG_TI_JMB_FRAMES   (0),
  .CFG_NSC_OPERATION   (0)
)USPIM ( //.TESTMODE   (1'b0),
                  .PCLK       (PCLK),   
                  .PRESETN    (PRESETN),
                  .PADDR      (PADDR[6:0]),  
                  .PSEL       (PSEL[0]),   
                  .PENABLE    (PENABLE),
                  .PWRITE     (PWRITE), 
                  .PWDATA     (PWDATA), 
                  .PRDATA     (PRDATA_0),

                  .SPISSI     (), 
                  .SPISDI     (S_SPISDO), 
                  .SPICLKI    (),
                  .SPISS      (M_SPISS),  
                  .SPISCLKO   (M_SPISCLKO),  
                  .SPIOEN     (M_SPIOEN),    
                  .SPISDO     (M_SPISDO),    

                  .SPIINT     (GP_IN[0]), 
                  .SPIRXAVAIL (),
                  .SPITXRFM   (),  
                  .SPIMODE    (),
                  .PREADY     (),
                  .PSLVERR    ()

                  );

// ********************************************************************************
// SPI Core - Slave  

wire [7:0] S_SPISS;


CORESPI # (
  //.FAMILY              (FAMILY),
  .APB_DWIDTH          (32),
  .CFG_FRAME_SIZE      (32),
  .CFG_FIFO_DEPTH      (4),
  .CFG_CLK             (3),
  .CFG_MODE            (0),
  .CFG_MOT_MODE        (0),
  .CFG_MOT_SSEL        (0),
  .CFG_TI_NSC_CUSTOM   (0),
  .CFG_TI_NSC_FRC      (0),
  .CFG_TI_JMB_FRAMES   (0),
  .CFG_NSC_OPERATION   (0)
)  USPIS ( //.TESTMODE   (1'b0),
                  .PCLK       (PCLK),   
                  .PRESETN    (PRESETN),
                  .PADDR      (PADDR[6:0]),  
                  .PSEL       (PSEL[1]),   
                  .PENABLE    (PENABLE),
                  .PWRITE     (PWRITE), 
                  .PWDATA     (PWDATA), 
                  .PRDATA    (PRDATA_1),

                  .SPISSI     (M_SPISS[0]), 
                  .SPISDI     (M_SPISDO), 
                  .SPICLKI    (M_SPISCLKO),
                  .SPISS      (),  
                  .SPISCLKO   (),  
                  .SPIOEN     (),    
                  .SPISDO     (S_SPISDO),    

                  .SPIINT     (GP_IN[1]), 
                  .SPIRXAVAIL (),
                  .SPITXRFM   (),  
                  .SPIMODE    (),
                  .PREADY     (),
                  .PSLVERR    ()
                  );
endmodule

